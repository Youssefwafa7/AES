module adder (in, out,outing);
    input in;
    output out,outing;
    assign out = in;
    assign outing = in;
endmodule