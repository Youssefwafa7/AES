module adder (in, out,og);
    input in;
    output out,og;
    assign out = in;
    assign og = in;
    //trying commits
endmodule