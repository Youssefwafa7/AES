module SubBytes(input [0:31] in , output [0:31] out);



endmodule