module Cipher (state_in , keys , state_out);
    input [127:0]state_in;
    input [1407:0]keys;  
    output [127:0]state_in;
    



endmodule